// Instruction type
`define R_TYPE 7'b0110011 //Register to Register(Arthmetic and Logical)
`define I_TYPE 7'b0010011 //Immediate Operations
`define S_TYPE 7'b0100011 //Store Instructions
`define B_TYPE 7'b1100011 //Branch Instructions
`define U_TYPE 7'b0110111 //Load Instructions
`define J_TYPE 7'b1101111 //Jump Instructions
