module instruction_tb;

 

endmodule
