// Instruction type
`define R_TYPE 7'b0110011 //Register to Register(Arthmetic and Logical)
`define I_TYPE 7'b0010011 //Immediate Operations
`define L_TYPE 7'b0000011 //Load Operations
`define S_TYPE 7'b0100011 //Store Instructions
`define B_TYPE 7'b1100011 //Branch Instructions
`define U_TYPE 7'b0110111 //Upper Immediate Instructions
`define J_TYPE 7'b1101111 //Jump Instructions
